module game (
    input wire pixel_clk_in,
    input wire rst_in,
    input wire start_btn,
    
    output logic game_state //TODO: SET BITS
    
)

endmodule