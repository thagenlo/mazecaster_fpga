`timescale 1ns / 1ps
`default_nettype none

module transformation

endmodule

`default_nettype wire