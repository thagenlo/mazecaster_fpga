// module game_fsm #(
//     parameter ROTATION_ANGLE = 16'b0010_1101_0000_0000 // default = 45 degrees
//     )(input wire clk_in,
//     input wire rst_in,
//     input wire [15:0] posX, 
//     input wire [15:0] posY,
//     output logic state 
//     );


// endmodule